`include "cpu_synth.v"
`include "memory.v"
`include "interruptcontroller.v"
`include "timer.v"
`include "gpio.v"
`include "watchdog.v"

`begin_keywords "1800-2009"

`timescale 1us/1ns

module clkgen (clk);
	output reg clk;

	initial
		clk = 0;

	always #5 clk = !clk;
endmodule

module iosystem
	#(parameter
	IRQCTRLADDRBASE = 16'h0010,
	TIMER0ADDRBASE = 16'h0018,
	WATCHDOGADDRBASE = 16'h0020,
	GPIO0ADDDRBASE = 16'h0028)
	
	(input logic [15:0] dread_addr, output logic [15:0] dread_data,
	input logic [15:0] dwrite_addr, dwrite_data, input logic [1:0] dwrite_en,
	output logic interrupt, input logic clk, output logic reset, input logic trap, input logic power_on_reset);

	wire [15:0] dwrite_addr_even, dwrite_addr_odd;
	wire [15:0] dread_addr_even, dread_addr_odd;
	wire dwrite_en_even, dwrite_en_odd;
	assign dread_addr_even = dread_addr[0] ? dread_addr + 1 : dread_addr;
	assign dread_addr_odd = dread_addr[0] ? dread_addr : dread_addr + 1;
	assign dwrite_addr_even = dwrite_addr[0] ? dwrite_addr + 1 : dwrite_addr;
	assign dwrite_addr_odd = dwrite_addr[0] ? dwrite_addr : dwrite_addr + 1;
	assign dwrite_en_even = dwrite_addr[0] ? dwrite_en[1] : dwrite_en[0];
	assign dwrite_en_odd = dwrite_addr[0] ? dwrite_en[0] : dwrite_en[1];

	// Interrupt controller
	wire irqctrl_enable_read, irqctrl_active_read;
	wire irqctrl_enable_write, irqctrl_active_write;
	wire timer_counter_write[1:0], timer_reload_write[1:0], timer_config_write;
	logic [1:0] irqctrl_enable_dread, irqctrl_active_dread;
	logic [1:0] irqctrl_enable_dwrite, irqctrl_active_dwrite;
	logic [1:0] interrupts;
	assign irqctrl_enable_read = (dread_addr_even == IRQCTRLADDRBASE);
	assign irqctrl_active_read = (dread_addr_even == IRQCTRLADDRBASE + 2);
	assign irqctrl_enable_write = dwrite_en_even && (dwrite_addr_even == IRQCTRLADDRBASE);
	assign irqctrl_active_write = dwrite_en_even && (dwrite_addr_even == IRQCTRLADDRBASE + 2);
	interruptcontroller #(.NUM_INPUTS(2))
		irqctrl(.int_out(interrupt), .enable_out(irqctrl_enable_dread), .active_out(irqctrl_active_dread), .enable_in(dwrite_data[1:0]), .active_in(dwrite_data[1:0]), .enable_in_write(irqctrl_enable_write), .active_in_write(irqctrl_active_write),
		.in(interrupts), .*);

	// Timer 0
	wire timer0ovirq, timer0cmpirq;
	logic [0:0] timer0in;
	logic [1:0] timer0_counter_write, timer0_reload_write, timer0_compare_write;
	logic timer0_config_read;
	logic timer0_config_write;
	logic [7:0] timer0_config_dread;
	logic [15:0] timer0_counter_dread, timer0_reload_dread, timer0_compare_dread;
	logic [7:0] timer0_config_dwrite;
	logic [15:0] timer0_counter_dwrite, timer0_reload_dwrite, timer0_compare_dwrite;
	assign interrupts[0] = timer0ovirq;
	assign interrupts[1] = timer0cmpirq;
	always_comb
	begin
		timer0_config_read = (dread_addr_even == TIMER0ADDRBASE);
		timer0_config_write = dwrite_en_even && (dwrite_addr_even == TIMER0ADDRBASE);
		timer0_counter_write = {dwrite_en_odd && (dwrite_addr_odd == TIMER0ADDRBASE + 3), dwrite_en_even && (dwrite_addr_even == TIMER0ADDRBASE + 2)};
		timer0_reload_write = {dwrite_en_odd && (dwrite_addr_odd == TIMER0ADDRBASE + 5), dwrite_en_even && (dwrite_addr_even == TIMER0ADDRBASE + 4)};
		timer0_compare_write = {dwrite_en_odd && (dwrite_addr_odd == TIMER0ADDRBASE + 7), dwrite_en_even && (dwrite_addr_even == TIMER0ADDRBASE + 6)};
	end
	timer timer0(.counter_out(timer0_counter_dread), .reload_out(timer0_reload_dread), .compare_out(timer0_compare_dread), .config_out(timer0_config_dread),
		.overflow_int(timer0ovirq), .compare_int(timer0cmpirq), .counter_in(dwrite_data), .reload_in(dwrite_data), .compare_in(dwrite_data), .config_in(dwrite_data[7:0]),
		.counter_write(timer0_counter_write), .reload_write(timer0_reload_write), .compare_write(timer0_compare_write), .config_write(timer0_config_write), .in(timer0in), .*);

	// Watchdog
	logic [1:0] watchdog_counter_write, watchdog_reload_write;
	logic watchdog_config_read;
	logic watchdog_config_write;
	logic [7:0] watchdog_config_dread;
	logic [15:0] watchdog_counter_dread, watchdog_reload_dread;
	logic [7:0] watchdog_config_dwrite;
	logic [15:0] watchdog_counter_dwrite, watchdog_reload_dwrite;
	always_comb
	begin
		watchdog_config_read = (dread_addr_even == WATCHDOGADDRBASE);
		watchdog_config_write = dwrite_en_even && (dwrite_addr_even == WATCHDOGADDRBASE);
		watchdog_counter_write = {dwrite_en_odd && (dwrite_addr_odd == WATCHDOGADDRBASE + 3), dwrite_en_even && (dwrite_addr_even == WATCHDOGADDRBASE + 2)};
		watchdog_reload_write = {dwrite_en_odd && (dwrite_addr_odd == WATCHDOGADDRBASE + 5), dwrite_en_even && (dwrite_addr_even == WATCHDOGADDRBASE + 4)};
	end
	watchdog watchdog(.counter_out(watchdog_counter_dread), .reload_out(watchdog_reload_dread), .config_out(watchdog_config_dread),
		.counter_in(dwrite_data), .reload_in(dwrite_data), .config_in(dwrite_data[7:0]),
		.counter_write(watchdog_counter_write), .reload_write(watchdog_reload_write), .config_write(watchdog_config_write), .*);

	always @(posedge clk)
	begin
		if (dread_addr_even == dwrite_addr_even)
			dread_data[7:0] = dwrite_data;
		else if (irqctrl_enable_read)
			dread_data[7:0] = {'x, irqctrl_enable_dread[0:0]};
		else if (irqctrl_active_read)
			dread_data[7:0] = {'x, irqctrl_active_dread[0:0]};
		else if (timer0_config_read)
			dread_data[7:0] = {'x, timer0_config_dread[7:0]};
		else
			dread_data[7:0] = 'x;
		if (dread_addr_odd == dwrite_addr_odd)
			dread_data[15:8] = dwrite_data;
		else
			dread_data[15:8] = 'x;
	end
endmodule

module testsystem ();
	parameter RAMADDRBASE = 16'h2000;
	
	wire [15:0] iread_addr, dread_addr, dwrite_addr;
	wire [23:0] iread_data;
	logic [15:0] dread_data, dwrite_data;
	wire iread_valid;
	wire [1:0] dwrite_en;
	wire clk;
	reg power_on_reset;
	wire reset;
	wire interrupt;
	wire trap;

	wire [1:0] mem_dwrite_en, io_dwrite_en;
	wire [15:0] mem_dread_data, io_dread_data;

	clkgen clkgen(.*);
	cpu cpu(.*);
	memory memory(.dwrite_en(mem_dwrite_en), .dread_data(mem_dread_data), .*);
	iosystem iosystem(.dwrite_en(io_dwrite_en), .dread_data(io_dread_data), .*);

	logic [15:0] old_dread_addr;
	always @(posedge clk)
	begin
		old_dread_addr = dread_addr;
	end

	assign mem_dwrite_en = (dwrite_addr >= RAMADDRBASE) ? dwrite_en : 2'b00;
	assign io_dwrite_en = (dwrite_addr < RAMADDRBASE) ? dwrite_en : 2'b00;

	always_comb
	begin
		if (old_dread_addr >= RAMADDRBASE)
			dread_data = mem_dread_data;
		else
			dread_data = io_dread_data;
	end

	initial
	begin
		$dumpfile("postsynthcputest.vcd");
    	$dumpvars(0,testsystem);
    	power_on_reset <= 1;
    	#20
    	power_on_reset <= 0;
		#2180
		$finish;
	end

	always @(posedge trap)
	begin
		$display("ERROR: TRAP");
		#20
		$finish;
	end
endmodule

`end_keywords

